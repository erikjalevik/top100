Poisecore feat. Hannah Stacia\Lost In The Music\2017\2018\1
DJ Seinfeld\Time Spent Away From U\2017\2018\2
Technikore & UFO feat. Scandal\Always\2011\2018\3
Kim Petras\I Don't Want It At All\2017\2018\4
John Maus\Drinking Song\2018\2018\5
Alice Coltrane\Journey to Satchidananda\2017\2018\6
Drab Majesty\Dot in the Sky\2017\2018\7
DJ Seinfeld\U\2017\2018\8
Nadja\Sunwell\2018\2018\9
Da Tweekaz\Hewwego (Darren Styles Remix)\2016\2018\10
Converge\All We Love We Leave Behind\2012\2018\11
Charli XCX feat. Hannah Diamond\Paradise\2016\2018\12
Kælan Mikla\Kalt (Live)\2016\2018\13
Hannah Diamond\Fade Away\2016\2018\14
Hannah Diamond\Hi\2016\2018\15
Hannah Diamond\Never Again\2017\2018\16
Caterina Barbieri\Gravity that Binds\2017\2018\17
Nouvelle Phénomène\Cruel Game (Vanzetti & Sacco Remix)\2015\2018\18
DJ Seinfeld\U Hold Me Without Touch\2017\2018\19
Nabihah Iqbal\Zone 1 to 6000\2017\2018\20
A. G. Cook\Superstar\2016\2018\21
K Rizz\Imagine If\2014\2018\22
DJ Seinfeld\Too Late For U And M1\2017\2018\23
John Maus\Dumpster Baby\2018\2018\24
Cold Cave\Glory\2017\2018\25
Alice Coltrane\Krishna Krishna\1982\2018\26
DJ Seinfeld\I Hope I Sleep Tonight\2017\2018\27
Caterina Barbieri\SOTRS\2017\2018\28
Teengirl Fantasy\Star-Rise\2017\2018\29
DJ Seinfeld\I Saw Her Kiss Him In Front Of Me And I Was Like Wtf?\2017\2018\30
Farah\Into Eternity (Main)\2013\2018\31
Null+Void feat. Dave Gahan\Where I Wait\2017\2018\32
Lords of Midnite\Drown in Ur Love\2013\2018\33
DJ DJ Booth\Heaven (A.G. Cook Remix)\2013\2018\34
Fraunhofer Diffraction\My Baby\2013\2018\35
Collapse\My Love (Ambient Drops)\1991\2018\36
Venetian Snares\Everything About You Is Special\2016\2018\37
DJ Seinfeld\Come Thru For U\2017\2018\38
Legowelt\Axumisia V S612\2017\2018\39
Marquis Hawkes feat. Ursula Rucker\Don't U (Edit)\2018\2018\40
CFCF\Cell Site in Somerset\2018\2018\41
Robyn\Because It's In The Music\2018\2018\42
Nightwish\Dark Chest of Wonders\2004\2018\43
Austra\American Science\2014\2018\44
Charli XCX feat. Kim Petras and Jay Park\Unlock It\2017\2018\45
Fraunhofer Diffraction\Kvrt In Space\2013\2018\46
Blonde feat. Alex Newell\All Cried Out\2015\2018\47
Babymetal\Megitsune\2014\2018\48
Giuseppe Ottaviani feat. Hypaton\Space Unicorn\2018\2018\49
Black Loops\Get Lost\2016\2018\50
Nadja\In The Shadow Of The Wing Of The Thing Too Big To Be Seen\2018\2018\51
Marquis Hawkes feat. Jocelyn Brown\I'm So Glad (Paul Woolford Rework)\2016\2018\52
John O'Callaghan feat. Josie\Out Of Nowhere (Giuseppe Ottaviani Extended Remix)\2018\2018\53
Trisomie 21\The Last Song\1986\2018\54
Alice Coltrane\Keshava Murahara\2017\2018\55
Jimmy Edgar feat. Dawn\Burn So Deep (Extended Mix)\2018\2018\56
Microwave Prince\Microwavin'\1993\2018\57
The Blaze\Territory\2017\2018\58
Reso\Kodama\2017\2018\59
DJ Q feat. Louise Williams\Through The Night (Deckstar Vocal 2step Mix)\2013\2018\60
Hannah Diamond\Make Believe\2016\2018\61
Giuseppe Ottaviani\Ozone (Craig Connelly Extended Remix)\2018\2018\62
Paul Van Dyk\My World (Florjn Mix)\1994\2018\63
Robyn\Send To Robin Immediately\2018\2018\64
Brisk & Vinylgroover\Checkin' Da Cutz (M-Project & Liqo Remix)\2017\2018\65
Tangerine Dream\Sensing Elements\2017\2018\66
ionnalee feat. Jamie Irrepressible\Dunes of Sand\2018\2018\67
Rebekah\Waiting For You\2018\2018\68
Caterina Barbieri\Scratches on the Readable Surface\2017\2018\69
Babymetal\Iine!\2014\2018\70
DJ Seinfeld\With My Luv\2017\2018\71
Imre Kiss\You And Me Are The Same\2018\2018\72
Rival Consoles\Untravel\2018\2018\73
Julee Cruise\Questions in a World of Blue\1993\2018\74
Tommy 86 feat. Sally Shapiro\Why Did I Say Goodbye\2014\2018\75
Popsimonova\Drive\2015\2018\76
Plus System\This Is How We Do It\2004\2018\77
Reso\Avenoir\2018\2018\78
Hannah Diamond\Concrete Angel\2017\2018\79
Both Hands Free\Phobos\1976\2018\80
Special Request\Brainstorm (Gerd Janson & Shan House Mix)\2018\2018\81
Kedr Livanskiy\Ariadna\2017\2018\82
Randy Crawford\Just To Keep You Satisfied\1979\2018\83
Mister Shifter\Dreada\2018\2018\84
John Maus\Touchdown\2017\2018\85
Marquis Hawkes & Jamie Lidell\We Should Be Free (Hawkes Dub)\2018\2018\86
Against All Logic\Some Kind Of Game\2018\2018\87
Julee Cruise\In My Other World\1993\2018\88
Objekt\Ganzfeld\2014\2018\89
Teengirl Fantasy feat. Khalif Jones\Seeds\2017\2018\90
Reso\Aural Animation\2018\2018\91
Nightwish\Ghost Love Score\2004\2018\92
Hercules & Love Affair Feat. John Grant\I Try To Talk To You\2014\2018\93
Kim Petras\In The Next Life\2018\2018\94
Black Ivory\Mainline\1979\2018\95
Kim Petras\Close Your Eyes\2018\2018\96
Robyn\Honey\2018\2018\97
Teengirl Fantasy\Crash Soft\2017\2018\98
Let's Eat Grandma\Hot Pink\2018\2018\99
Jakka-B\Lost In The Rhythm\2017\2018\100
