2016\1\AU
2016\1\UK
2016\2\DE
2016\3\NO
2016\4\US
2016\5\UK
2016\6\UK
2016\7\UK
2016\8\UK
2016\9\UK
2016\10\UK
2016\11\NL
2016\12\UK
2016\13\UK
2016\14\IT
2016\15\DE
2016\16\UK
2016\17\AU
2016\17\UK
2016\18\US
2016\19\UK
2016\20\US
2016\21\SE
2016\22\UK
2016\23\UK
2016\24\UK
2016\25\UK
2016\26\UK
2016\27\UK
2016\28\UK
2016\29\UK
2016\30\UK
2016\31\DE
2016\32\IT
2016\33\US
2016\34\DE
2016\35\AU
2016\35\UK
2016\36\US
2016\37\US
2016\38\UK
2016\39\DE
2016\39\UA
2016\40\UK
2016\41\UK
2016\42\NG
2016\43\UK
2016\44\AU
2016\44\UK
2016\45\UK
2016\46\DE
2016\47\UK
2016\48\NL
2016\49\UK
2016\50\UK
2016\51\US
2016\52\UK
2016\53\UK
2016\54\NO
2016\54\UK
2016\55\UK
2016\56\KW
2016\57\ES
2016\58\UK
2016\59\JP
2016\60\UK
2016\61\UK
2016\62\US
2016\63\UK
2016\64\US
2016\65\UK
2016\66\NG
2016\67\UK
2016\68\CA
2016\68\US
2016\69\KW
2016\70\UK
2016\71\NL
2016\71\UA
2016\72\UK
2016\73\UK
2016\74\UK
2016\75\US
2016\75\DE
2016\76\UK
2016\77\UK
2016\78\US
2016\79\UK
2016\80\NO
2016\81\DE
2016\82\UK
2016\83\VE
2016\84\DE
2016\85\US
2016\86\DE
2016\86\UK
2016\87\UK
2016\88\UK
2016\89\US
2016\89\DE
2016\90\UK
2016\91\US
2016\92\UK
2016\93\US
2016\94\UK
2016\95\US
2016\96\UK
2016\97\UK
2016\98\FI
2016\99\UK
2016\100\UK
2014\1\UK
2014\2\UK
2014\3\UK
2014\4\UK
2014\5\UK
2014\6\UK
2014\7\UK
2014\8\UK
2014\9\UK
2014\10\UK
2014\11\UK
2014\12\NL
2014\13\DE
2014\13\UK
2014\14\CA
2014\14\US
2014\15\UK
2014\16\UK
2014\17\UK
2014\17\FR
2014\18\UK
2014\19\NL
2014\20\UK
2014\21\DE
2014\22\UK
2014\23\US
2014\24\UK
2014\25\US
2014\26\DE
2014\27\UK
2014\28\US
2014\29\UK
2014\30\US
2014\31\UK
2014\32\UK
2014\33\NL
2014\34\US
2014\35\US
2014\36\US
2014\37\RU
2014\38\UK
2014\39\DE
2014\40\FR
2014\41\SE
2014\42\US
2014\43\FR
2014\43\US
2014\44\UK
2014\45\UK
2014\46\US
2014\47\US
2014\48\UK
2014\49\UK
2014\50\UK
2014\51\DE
2014\52\US
2014\53\IE
2014\53\IT
2014\54\UK
2014\55\IT
2014\56\US
2014\57\LT
2014\58\UK
2014\59\UK
2014\60\ES
2014\61\UK
2014\62\UK
2014\63\US
2014\64\UK
2014\65\FR
2014\66\UK
2014\67\UK
2014\68\UK
2014\69\SE
2014\69\NL
2014\70\UK
2014\71\UK
2014\72\UK
2014\73\US
2014\74\DE
2014\75\US
2014\76\DE
2014\77\DE
2014\78\DE
2014\79\DE
2014\80\US
2014\81\JP
2014\82\US
2014\83\UK
2014\84\CA
2014\85\UK
2014\86\US
2014\87\RU
2014\88\RU
2014\89\UK
2014\90\UK
2014\91\UK
2014\92\US
2014\93\RU
2014\94\UK
2014\95\UK
2014\96\UK
2014\97\UK
2014\98\US
2014\99\IT
2014\100\DE
2013\1\CA
2013\2\ZA
2013\2\UK
2013\3\UK
2013\4\UK
2013\5\UK
2013\6\SE
2013\7\UK
2013\8\US
2013\9\NL
2013\10\UK
2013\11\SE
2013\12\UK
2013\13\UK
2013\14\US
2013\15\US
2013\16\US
2013\17\US
2013\18\US
2013\19\US
2013\20\SE
2013\21\DE
2013\22\FR
2013\23\DK
2013\23\UK
2013\24\US
2013\25\US
2013\26\UK
2013\27\UK
2013\28\UK
2013\29\US
2013\30\US
2013\31\HU
2013\32\UK
2013\33\US
2013\34\UK
2013\35\SE
2013\36\IT
2013\37\US
2013\38\CA
2013\39\SE
2013\40\US
2013\41\ES
2013\42\UK
2013\43\US
2013\44\US
2013\45\UK
2013\46\UK
2013\47\US
2013\48\SE
2013\49\UK
2013\50\US
2013\51\UK
2013\52\US
2013\53\SE
2013\54\UK
2013\55\ZA
2013\56\SE
2013\57\NL
2013\58\UK
2013\59\US
2013\60\SE
2013\61\UK
2013\62\UK
2013\63\CA
2013\64\NO
2013\65\SE
2013\66\DE
2013\67\UK
2013\68\UK
2013\69\LB
2013\70\SE
2013\71\DE
2013\72\NO
2013\73\US
2013\74\US
2013\75\DE
2013\76\BE
2013\77\SE
2013\78\UK
2013\79\UK
2013\80\UK
2013\81\UK
2013\82\UK
2013\83\FR
2013\84\US
2013\85\UK
2013\86\UK
2013\87\UK
2013\88\US
2013\88\UK
2013\89\IN
2013\90\US
2013\91\UK
2013\92\UK
2013\93\UK
2013\94\SE
2013\95\NO
2013\96\US
2013\97\US
2013\98\US
2013\99\UK
2013\100\UK
2012\1\US
2012\2\US
2012\3\US
2012\3\UK
2012\4\US
2012\5\US
2012\6\DE
2012\7\UK
2012\8\CA
2012\9\UK
2012\10\US
2012\11\GE
2012\12\UK
2012\13\DE
2012\14\US
2012\15\UK
2012\16\UK
2012\17\DE
2012\18\UK
2012\19\UK
2012\20\US
2012\21\SE
2012\22\DE
2012\23\UK
2012\24\UK
2012\25\UK
2012\26\IS
2012\26\DE
2012\27\US
2012\28\IT
2012\29\UK
2012\30\DE
2012\30\FR
2012\31\CA
2012\32\IT
2012\33\FR
2012\33\CA
2012\34\US
2012\35\SE
2012\36\ES
2012\37\CA
2012\38\US
2012\39\NO
2012\40\US
2012\41\CA
2012\42\UK
2012\42\US
2012\43\US
2012\44\UK
2012\45\UK
2012\46\DE
2012\46\UA
2012\47\UK
2012\48\NL
2012\49\UK
2012\50\FI
2012\51\UK
2012\52\US
2012\53\UK
2012\54\IS
2012\54\DE
2012\55\HU
2012\56\UK
2012\57\UK
2012\58\UK
2012\59\US
2012\60\UK
2012\61\CA
2012\62\US
2012\63\UK
2012\64\CA
2012\64\US
2012\65\ES
2012\66\US
2012\67\UK
2012\68\UK
2012\69\LV
2012\70\DE
2012\71\DE
2012\72\US
2012\73\UK
2012\74\UK
2012\75\CA
2012\76\UK
2012\76\DE
2012\77\US
2012\78\NL
2012\79\CA
2012\80\IN
2012\81\UK
2012\82\ES
2012\83\US
2012\84\US
2012\85\FR
2012\86\US
2012\87\UK
2012\88\UK
2012\89\NZ
2012\89\UK
2012\90\CA
2012\91\IT
2012\92\FR
2012\93\NL
2012\94\US
2012\95\UK
2012\96\US
2012\97\DE
2012\98\US
2012\99\UK
2012\100\SE
2011\1\UK
2011\2\ES
2011\3\US
2011\4\US
2011\5\FR
2011\6\US
2011\7\SE
2011\8\UK
2011\9\IT
2011\10\US
2011\11\US
2011\12\NO
2011\13\UK
2011\14\UK
2011\15\US
2011\16\UK
2011\17\UK
2011\18\UK
2011\19\UK
2011\20\DE
2011\21\FR
2011\21\NL
2011\22\US
2011\23\CA
2011\24\DE
2011\25\NO
2011\26\US
2011\27\CA
2011\28\US
2011\29\SE
2011\30\FR
2011\31\US
2011\32\US
2011\33\UK
2011\34\NO
2011\35\US
2011\36\ES
2011\37\NL
2011\38\US
2011\39\FI
2011\40\US
2011\41\UK
2011\42\US
2011\43\US
2011\43\CA
2011\44\US
2011\45\CA
2011\46\DE
2011\47\IT
2011\48\UA
2011\48\DE
2011\49\US
2011\50\NO
2011\51\US
2011\52\UK
2011\53\UK
2011\54\SE
2011\55\NO
2011\56\UK
2011\57\US
2011\58\US
2011\59\IT
2011\60\UK
2011\61\US
2011\62\UK
2011\63\US
2011\63\DE
2011\64\UK
2011\65\CA
2011\66\SE
2011\67\US
2011\68\US
2011\69\NL
2011\70\UK
2011\71\NL
2011\72\SE
2011\73\SE
2011\74\IT
2011\75\CA
2011\76\DE
2011\77\FR
2011\78\US
2011\79\CA
2011\80\SE
2011\81\US
2011\82\ES
2011\83\IT
2011\84\UK
2011\85\UK
2011\86\US
2011\87\US
2011\88\UK
2011\89\UK
2011\90\NZ
2011\91\SE
2011\92\LV
2011\93\US
2011\94\UK
2011\95\NO
2011\96\AT
2011\96\SE
2011\97\UK
2011\98\UK
2011\99\DE
2011\100\UK
2010\1\US
2010\2\US
2010\3\US
2010\4\US
2010\5\US
2010\6\US
2010\7\US
2010\8\AR
2010\9\UK
2010\10\US
2010\11\US
2010\12\US
2010\12\CA
2010\13\SE
2010\14\US
2010\15\US
2010\16\US
2010\17\AT
2010\18\US
2010\19\DE
2010\20\US
2010\21\UK
2010\22\US
2010\23\US
2010\24\US
2010\25\US
2010\26\US
2010\27\US
2010\28\IT
2010\29\FR
2010\30\US
2010\31\US
2010\32\US
2010\33\US
2010\34\UK
2010\35\US
2010\36\SE
2010\37\US
2010\38\US
2010\39\UK
2010\40\IT
2010\41\RS
2010\42\US
2010\43\DE
2010\44\US
2010\45\SE
2010\46\US
2010\47\US
2010\48\FI
2010\49\CA
2010\49\US
2010\50\US
2010\51\UK
2010\52\UK
2010\53\US
2010\54\UK
2010\55\US
2010\56\US
2010\57\US
2010\58\US
2010\59\US
2010\60\BE
2010\61\US
2010\62\US
2010\63\US
2010\64\UK
2010\65\US
2010\66\US
2010\67\IT
2010\67\US
2010\68\CA
2010\69\SE
2010\70\US
2010\71\US
2010\72\IT
2010\73\SE
2010\74\SE
2010\75\DE
2010\76\UK
2010\77\DE
2010\78\US
2010\79\US
2010\80\SE
2010\81\FR
2010\82\UK
2010\83\IT
2010\84\US
2010\85\US
2010\86\US
2010\87\SE
2010\88\NL
2010\89\US
2010\90\SE
2010\91\IT
2010\92\US
2010\93\DE
2010\94\US
2010\95\US
2010\96\US
2010\97\UK
2010\98\US
2010\99\CA
2010\100\UK
2009\1\IT
2009\2\DE
2009\2\US
2009\3\DE
2009\3\US
2009\4\FR
2009\5\US
2009\6\US
2009\7\IL
2009\8\DE
2009\9\US
2009\10\ZA
2009\11\SE
2009\12\FI
2009\13\US
2009\13\UK
2009\14\DE
2009\15\UK
2009\16\SE
2009\17\US
2009\18\FR
2009\19\ES
2009\20\US
2009\21\SE
2009\22\NL
2009\23\UK
2009\24\SE
2009\25\SE
2009\26\UK
2009\27\US
2009\28\SE
2009\29\FR
2009\30\US
2009\30\CA
2009\31\NL
2009\32\US
2009\33\UK
2009\34\UK
2009\35\US
2009\36\US
2009\37\UK
2009\37\US
2009\37\IT
2009\37\BE
2009\38\NO
2009\39\UK
2009\40\UK
2009\41\DE
2009\41\US
2009\42\DE
2009\43\IT
2009\44\IT
2009\45\UK
2009\46\US
2009\47\US
2009\48\DE
2009\49\SE
2009\50\NL
2009\51\US
2009\51\UK
2009\52\US
2009\53\NL
2009\54\US
2009\55\DE
2009\56\US
2009\57\UK
2009\58\DE
2009\59\SE
2009\60\US
2009\61\FI
2009\62\SE
2009\63\US
2009\64\UK
2009\65\UK
2009\66\US
2009\67\CA
2009\68\FI
2009\69\SE
2009\70\US
2009\71\UK
2009\72\UK
2009\73\UK
2009\74\UK
2009\75\US
2009\76\UK
2009\77\AU
2009\77\US
2009\78\US
2009\79\FI
2009\80\IT
2009\80\BE
2009\81\UK
2009\82\US
2009\83\NL
2009\84\CA
2009\85\US
2009\85\NL
2009\86\UK
2009\87\IT
2009\88\NL
2009\89\US
2009\90\UK
2009\91\ES
2009\91\NL
2009\92\NL
2009\93\UK
2009\94\CA
2009\94\US
2009\95\UK
2009\96\UK
2009\97\SE
2009\98\UK
2009\99\FR
2009\100\US
2008\1\SE
2008\2\US
2008\3\SE
2008\4\DE
2008\4\FR
2008\5\SE
2008\6\SE
2008\7\DE
2008\8\SE
2008\9\US
2008\10\SE
2008\11\FR
2008\12\US
2008\13\US
2008\14\CA
2008\15\PL
2008\16\NL
2008\17\PL
2008\18\DE
2008\19\UK
2008\20\UK
2008\21\SE
2008\22\NL
2008\23\UK
2008\24\SE
2008\25\SE
2008\26\US
2008\27\SE
2008\28\IT
2008\29\US
2008\30\IT
2008\31\NO
2008\32\NL
2008\32\FR
2008\33\UK
2008\34\NO
2008\35\NL
2008\36\US
2008\37\SE
2008\38\NL
2008\39\IT
2008\40\DE
2008\41\DE
2008\42\IT
2008\43\SE
2008\43\FR
2008\44\US
2008\45\DE
2008\46\NO
2008\47\US
2008\48\US
2008\49\DE
2008\50\SE
2007\1\IT
2007\2\NL
2007\3\SE
2007\4\NL
2007\5\SE
2007\6\US
2007\7\IT
2007\8\FR
2007\9\NL
2007\10\SE
2007\11\UK
2007\12\UK
2007\13\DE
2007\14\SE
2007\15\IT
2007\16\IT
2007\17\SE
2007\18\SE
2007\19\NL
2007\20\DE
2007\21\SE
2007\22\IT
2007\23\SE
2007\23\FR
2007\24\DE
2007\25\US
2007\26\UK
2007\27\FR
2007\28\SE
2007\29\IT
2007\30\IT
2007\31\IT
2007\32\UK
2007\33\SE
2007\34\FR
2007\35\IT
2007\36\NO
2007\37\IT
2007\37\NL
2007\38\UK
2007\39\JP
2007\40\IT
2007\41\SE
2007\42\UK
2007\42\US
2007\43\IT
2007\44\US
2007\45\DE
2007\46\US
2007\47\UK
2007\48\IT
2007\49\SE
2007\50\NL
2007\51\IT
2007\52\SE
2007\53\UK
2007\54\US
2007\55\SE
2007\56\IT
2007\57\DE
2007\58\PL
2007\59\FR
2007\60\US
2007\61\FR
2007\61\UK
2007\62\US
2007\63\IT
2007\64\FR
2007\65\SE
2007\66\DE
2007\67\UK
2007\68\NL
2007\69\IT
2007\70\IT
2007\71\FR
2007\72\SE
2007\73\US
2007\74\NL
2007\75\SE
2007\76\UK
2007\77\DE
2007\78\US
2007\79\ES
2007\80\UK
2007\81\IT
2007\82\UK
2007\83\SE
2007\84\UK
2007\85\UK
2007\86\UK
2007\87\IT
2007\88\BE
2007\88\FR
2007\89\FR
2007\90\NL
2007\91\US
2007\92\UK
2007\93\IT
2007\94\SE
2007\95\ES
2007\96\US
2007\97\US
2007\98\SE
2007\99\DE
2007\99\UK
2007\100\PL
2006\1\IT
2006\2\SE
2006\3\SE
2006\4\IT
2006\5\IT
2006\6\IT
2006\7\SE
2006\8\IT
2006\9\AU
2006\10\SE
2006\11\IT
2006\12\AT
2006\13\NL
2006\14\NL
2006\15\FI
2006\16\US
2006\17\UK
2006\18\US
2006\19\SE
2006\20\NL
2006\21\IT
2006\22\SE
2006\23\SE
2006\24\NL
2006\25\SE
2006\26\UK
2006\27\IE
2006\28\UK
2006\29\SE
2006\30\IT
2006\31\DK
2006\32\CN
2006\32\FR
2006\32\NL
2006\33\NL
2006\34\IT
2006\35\IE
2006\36\IT
2006\37\FR
2006\38\CA
2006\39\NL
2006\40\SE
2006\41\IT
2006\42\NL
2006\43\SE
2006\44\JP
2006\45\UK
2006\46\IT
2006\47\SE
2006\48\PL
2006\49\UK
2006\50\NL
2005\1\IT
2005\2\AU
2005\3\SE
2005\4\NL
2005\5\US
2005\6\UK
2005\7\SE
2005\8\FI
2005\9\FR
2005\10\SE
2005\11\FR
2005\12\SE
2005\12\AU
2005\13\UK
2005\14\CA
2005\15\IE
2005\16\UK
2005\17\IE
2005\18\UK
2005\19\UK
2005\20\UK
2005\21\NL
2005\22\DE
2005\23\UK
2005\24\NL
2005\25\UK
2005\26\IE
2005\27\NL
2005\28\SE
2005\29\US
2005\30\US
2005\31\UK
2005\32\UK
2005\33\RU
2005\34\NL
2005\35\SE
2005\36\UK
2005\37\SE
2005\38\SE
2005\39\UK
2005\40\NL
2005\41\US
2005\41\UK
2005\42\SE
2005\42\DK
2005\43\UK
2005\44\DK
2005\45\DE
2005\46\US
2005\46\UK
2005\47\SE
2005\48\UK
2005\48\DE
2005\49\CA
2005\50\CA
