2018\1\UK
2018\2\SE
2018\3\UK
2018\4\US
2018\4\DE
2018\5\US
2018\6\US
2018\7\US
2018\8\SE
2018\9\CA
2018\10\NO
2018\10\UK
2018\11\US
2018\12\UK
2018\13\IS
2018\14\UK
2018\15\UK
2018\16\UK
2018\17\IT
2018\18\HU
2018\19\SE
2018\20\UK
2018\21\UK
2018\22\PH
2018\23\SE
2018\24\US
2018\25\US
2018\26\US
2018\27\SE
2018\28\IT
2018\29\US
2018\30\SE
2018\31\US
2018\32\US
2018\32\UK
2018\33\NL
2018\34\UK
2018\35\RU
2018\36\UK
2018\37\CA
2018\38\SE
2018\39\NL
2018\40\UK
2018\40\US
2018\41\CA
2018\42\SE
2018\43\FI
2018\44\US
2018\45\UK
2018\45\US
2018\45\DE
2018\45\KR
2018\46\RU
2018\47\UK
2018\47\US
2018\48\JP
2018\49\IT
2018\50\IT
2018\51\CA
2018\52\UK
2018\52\US
2018\53\IE
2018\53\US
2018\53\IT
2018\54\FR
2018\55\US
2018\56\US
2018\57\DE
2018\58\FR
2018\59\UK
2018\60\UK
2018\61\UK
2018\62\IT
2018\62\UK
2018\63\DE
2018\64\SE
2018\65\UK
2018\66\DE
2018\67\SE
2018\67\UK
2018\68\UK
2018\69\IT
2018\70\JP
2018\71\SE
2018\72\HU
2018\73\UK
2018\74\US
2018\75\FR
2018\75\SE
2018\76\HR
2018\77\UK
2018\78\UK
2018\79\UK
2018\80\UK
2018\81\UK
2018\81\DE
2018\82\RU
2018\83\US
2018\84\US
2018\85\US
2018\86\UK
2018\87\CL
2018\87\US
2018\88\US
2018\89\UK
2018\90\US
2018\91\UK
2018\92\FI
2018\93\US
2018\94\US
2018\94\DE
2018\95\US
2018\96\US
2018\96\DE
2018\97\SE
2018\98\US
2018\99\UK
2018\100\UK
