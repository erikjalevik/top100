Dead Can Dance\Persephone (The Gathering of Flowers)\1987\2016\1
EQD\005B\2011\2016\2
Susanne Sundfør\Slowly\2015\2016\3
Martial Canterel\Teano\2014\2016\4
Royal-T feat. P Money\Cruel to be Kind\2012\2016\5
George FitzGerald feat. Boxed In\Full Circle\2015\2016\6
DJ Q feat. MC Bonez\You Wot (Club Mix)\2007\2016\7
Après\Chicago (Club Edit)\2015\2016\8
High Contrast & Clare Maguire\Who's Loving You (Part 2)\2014\2016\9
Shadow Child & Ben Pearce feat. Laurel\Nothing Ever Hurts\2015\2016\10
Noisecontrollers\Break the Show\2012\2016\11
Special Request\Amnesia\2015\2016\12
Zomby\SURF I\2015\2016\13
Donato Dozzy\Gol\2006\2016\14
The Panacea\Found a Lover\2004\2016\15
Billon\Slave to the Vibe\2015\2016\16
Dead Can Dance\Summoning of The Muse\1987\2016\17
Martial Canterel\Bulvár\2014\2016\18
Paul Woolford\MDMA\2015\2016\19
Terrence Parker feat. Merachka\Open Up Your Spirit\2014\2016\20
Johan Agebjörn, Le Prix & Lake Heartbeat\Watch The World Go By\2011\2016\21
Danny L. Harle\Forever\2015\2016\22
Hannah Diamond\Every Night\2015\2016\23
P Money\War Dub (Reply to Ghetts)\2010\2016\24
Equinox\Killa Sound (B-Key Remix)\2011\2016\25
The Squire of Gothos\Walkin Manz Klub\2013\2016\26
DJ S.K.T feat. Rae\Take Me Away\2015\2016\27
Special Request\Simulation\2015\2016\28
Bicep\Closing Sequence\2015\2016\29
easyFun\Laplander\2015\2016\30
Juliane Werding\Großstadtlichter (Kinky Lovers Edit)\1980\2016\31
East Wall\Ice of Fire\1991\2016\32
Void Vision\Hidden Hand\2014\2016\33
Heaven Shall Burn\Whatever it May Take\2002\2016\34
Jagwar Ma\Uncertainty (Mssingno Remix)\2014\2016\35
Slava\Girl Like Me\2013\2016\36
Deniece Williams\Free\1976\2016\37
µ-Ziq\Forger\2015\2016\38
The Panacea feat. Goldberg Variations & Untergang\Ryse & Shiiine\2014\2016\39
Kayper\4 Fingers\2015\2016\40
µ-Ziq\Monj2\2015\2016\41
William Onyeabor\Good Name\1983\2016\42
Sophie\Just Like We Never Said Goodbye\2015\2016\43
Dead Can Dance\Dawn of the Iconoclast\1987\2016\44
Shadow Child & Doorly\Climbin' (Piano Weapon)\2014\2016\45
Heaven Shall Burn\Implore the Darken Sky\2002\2016\46
Unicorn Kid\Need U\2012\2016\47
Noisecontrollers\Sludge\2012\2016\48
DJ Q\They Haven't Got a Chance\2012\2016\49
Zomby\Float\2008\2016\50
Pictureplane\Esoterrorist\2015\2016\51
Zomby\Euphoria\2008\2016\52
µ-Ziq\Ritm\2015\2016\53
Jenny Hval\Kingsize (Kelly Lee Owens Rework)\2016\2016\54
Zomby\We Got the Sound\2008\2016\55
Fatima Al Qadiri\Szechuan\2014\2016\56
Pional\It's All Over\2014\2016\57
Kuedo\In Your Sleep\2016\2016\58
Babymetal\Gimme Chocolate!!\2014\2016\59
Zomby\Where Were U in '92\2008\2016\60
Special Request\Reset it\2015\2016\61
Martial Canterel\Baltic Coast\2014\2016\62
Palms Trax\Sumo Acid Crew\2015\2016\63
Terrence Parker\The Back 9\2014\2016\64
µ-Ziq\Smeester\2015\2016\65
William Onyeabor\When the Going is Smooth & Good\1985\2016\66
Special Request\Undead\2013\2016\67
Junior Boys\Big Black Coat (Robert Hood Remix)\2016\2016\68
Fatima Al Qadiri\Shanghai Freeway\2014\2016\69
Konx-Om-Pax\Rainbow Bounce\2016\2016\70
The Hard Way\Pentagram of Coke\2013\2016\71
Citizen\So Submissive\2013\2016\72
Floating Points\Kuiper\2016\2016\73
Burial\Temple Sleeper\2015\2016\74
Juan Atkins & Moritz von Oswald present Borderland\Zeolites\2016\2016\75
Special Request\Soundboy Killer\2013\2016\76
Unicorn Kid\Chrome Lion\2011\2016\77
Void Vision\Sour\2014\2016\78
Deadboy\Return\2014\2016\79
Jaga Jazzist\Oban (Todd Terje Remix)\2015\2016\80
Pantha du Prince\Dream Yourself Awake\2016\2016\81
µ-Ziq\Taxi Sadness\2015\2016\82
Arca\Mutant\2016\2016\83
Shed\Leave Things\2010\2016\84
Martial Canterel\Gyors-Lassú\2014\2016\85
Westbam feat. Richard Butler\You Need the Drugs (Extended Version)\2013\2016\86
Special Request\Deranged\2013\2016\87
Tessela\Hackney Parrot (Special Request VIP)\2013\2016\88
Juan Atkins & Moritz von Oswald present Borderland\Riod\2016\2016\89
Kuedo\Slow Knife\2016\2016\90
Martial Canterel\And I Thought\2014\2016\91
Special Request\Vapour\2013\2016\92
Terrence Parker feat. Coco Street\Hiding In Your Love\2014\2016\93
Palms Trax\People of Tusk\2015\2016\94
Matrixxman\Case Closed\2013\2016\95
Marquis Hawkes\Tunnel\2014\2016\96
Kuedo\Hourglass\2016\2016\97
Jaakko Eino Kalevi\Deeper Shadows\2015\2016\98
George FitzGerald feat. Lawrence Hart\Call it Love (If You Want to)\2015\2016\99
New Order\Tutti Frutti\2015\2016\100
Real Lies\North Circular\2014\2014\1
Sophie\Nothing More to Say\2012\2014\2
Mssingno\XE2\2013\2014\3
Hannah Diamond\Attachment\2014\2014\4
Flava D\Home\2013\2014\5
Mosca\Bax\2011\2014\6
Flava D\Hold On\2013\2014\7
Warrior One\Only You\2014\2014\8
Bicep\Keep Keep\2012\2014\9
Hannah Wants\Over\2012\2014\10
Danny L. Harle\Broken Flowers\2013\2014\11
Lenzman\Empty Promise\2013\2014\12
Technical Itch vs. The Panacea\Semisation 2013\2013\2014\13
Tim Hecker & Daniel Lopatin\Vaccination (for Thomas Mann)\2012\2014\14
A. G. Cook\Beautiful\2014\2014\15
Royal-T & Flava D\On My Mind (Version One)\2014\2014\16
Sophie\Bipp (Tielsie Remix)\2013\2014\17
Mssingno\XE3\2013\2014\18
Lenzman\Broken Dreams (Makoto Remix)\2013\2014\19
Vince Watson\Magma\2014\2014\20
Current Value\Dark Rain\2006\2014\21
Linea Aspera\Malarone\2012\2014\22
Xeno & Oaklander\Lastly\2014\2014\23
Disclosure feat. London Grammar\Help Me Lose My Mind (Paul Woolford Remix)\2013\2014\24
Xeno & Oaklander\G. Bruno\2014\2014\25
Anthony Rother\Technokultur\2014\2014\26
George FitzGerald\I can Tell (by the Way You Move)\2013\2014\27
Terrence Parker\Saved Forever\2014\2014\28
Vince Watson\A Very Different World\2009\2014\29
Floorplan\Never Grow Old\2013\2014\30
Depeche Mode\All That's Mine\2013\2014\31
Claude Speeed\Ssoon\2012\2014\32
Alden Tyrell\Somehouse\2013\2014\33
Joey Anderson\Above the Cherry Moon\2013\2014\34
Oneohtrix Point Never\Chrome Country\2013\2014\35
Xeno & Oaklander\Nuage d'Ivoire\2014\2014\36
Unquote feat. Grimm\Paint My Wings\2011\2014\37
Vince Watson\Otherworldy\2009\2014\38
Anthony Rother\Automat\2014\2014\39
Le Matin\Very Best of Myself\2014\2014\40
Cliff Lothar\Running Out of Time\2013\2014\41
DJ Rashad\Rollin'\2013\2014\42
Tielsie\Hueboy (DJ Clap Remix)\2014\2014\43
Vince Watson\Aurelon 10\2014\2014\44
Citizen\As One\2014\2014\45
Color War\SOS (DJ Clap Remix)\2014\2014\46
Terekke\Bank 3\2013\2014\47
Technimatic\Intersection\2013\2014\48
Bicep\Stash\2013\2014\49
Vince Watson\Free Yourself\2014\2014\50
Current Value\The Edge Of The Cliff\2006\2014\51
DJ Roc\One Blood\2010\2014\52
Mano Le Tough\Primative People (Tale of Us Remix)\2013\2014\53
Linea Aspera\Lamanai\2012\2014\54
Lory D\B1 Untitled\2001\2014\55
Xeno & Oaklander\Jasmine Nights\2014\2014\56
Ten Walls\Gotham\2013\2014\57
Roly Porter\Cloud\2013\2014\58
Bicep & Ejeca\You\2012\2014\59
Blanc 1\It's All Over\2013\2014\60
Citizen\U Don't Know\2014\2014\61
Hannah Wants & Chris Lorenzo\Girls\2014\2014\62
Omar S\Rewind\2013\2014\63
Bicep\Snack Bar\2013\2014\64
Tielsie\Palette\2014\2014\65
Linea Aspera\Fer-De-Lance\2012\2014\66
Life Sim\Caladhort\2014\2014\67
Linea Aspera\Eviction\2012\2014\68
Pagan Sector\The Corpse Fell into the Hourglass\2014\2014\69
Thy Slaughter\Bronze\2014\2014\70
Burial\Hiders\2013\2014\71
Bicep & Omar Odyssey\Don't\2012\2014\72
Greg Beato\Dreamin\2013\2014\73
Acasual\Spring Theory\2013\2014\74
Greg Beato\Who's the Licho in Charge Ovaa Here\2013\2014\75
Anthony Rother\In Digital Dominus\2014\2014\76
Anthony Rother\Widerstand\2014\2014\77
Anthony Rother\Schöpfer\2014\2014\78
Anthony Rother\Netzwerk\2014\2014\79
Matrixxman\Venetian Mask\2014\2014\80
Perfume\Night Flight\2009\2014\81
Oneohtrix Point Never\Along\2013\2014\82
Linea Aspera\Synapse\2012\2014\83
Kallisti\Arc of Fire\2013\2014\84
Warrior One\NYC\2014\2014\85
DJ Rashad & Gant-Man\Heaven Sent\2011\2014\86
Unquote feat. Grimm\Memories Fade Away\2011\2014\87
Unquote\Hide Your Tears Because We are in Heaven\2011\2014\88
Bicep\The Game\2013\2014\89
Bicep\Courtside Drama\2013\2014\90
A. G. Cook\Close Your Eyes\2013\2014\91
Oneohtrix Point Never\Still Life\2013\2014\92
Unquote\Reverberation Box\2011\2014\93
Hot Since 82\Knee Deep in Louise (Shadow Child Remix)\2012\2014\94
A. G. Cook feat. Hannah Diamond\Keri Baby\2014\2014\95
Bicep\Satisfy\2013\2014\96
Royal-T & Flava D\On My Mind (Version Three)\2014\2014\97
Fred P\Emotive Vibrations\2012\2014\98
Visonia\Impossible Romance\2014\2014\99
Anthony Rother\Ich Bin Ewig\2014\2014\100
Trust\Gloryhole\2012\2013\1
Red 7\I Lost My Shoes on Acid\2013\2013\2
Om Unit\Ulysses (Reso's Different Drum Remix)\2012\2013\3
Steve feat. Patricia Edwards\Love Dynasty\2013\2013\4
Chvrches\Recover (Curxes' 1996 Remix)\2013\2013\5
Sally Shapiro\Architectured Love\2013\2013\6
Photodementia\Refractivation\2013\2013\7
DJ Clap\Find Me a Lover\2011\2013\8
I-F\Superman (Live at the Bruine Planeet)\1995\2013\9
Disclosure feat. AlunaGeorge\White Noise\2013\2013\10
Sally Shapiro\If it doesn't Rain\2013\2013\11
Ital Tek\Yesterday Tomorrow Today\2012\2013\12
Disclosure feat. Sasha Keable\Voices\2013\2013\13
3 Channels\I can Understand\2011\2013\14
Black Marble\Pretender\2012\2013\15
Light Asylum\Hour Fortress\2012\2013\16
Underground Solution\Luv Dancin'\1990\2013\17
Light Asylum\Dark Allies\2010\2013\18
DJ Clap\Come On\2011\2013\19
Sally Shapiro\I Dream with an Angel Tonight\2013\2013\20
Die Selektion\Faust\2013\2013\21
Wax\Wax Dance (Dupe Edit)\1984\2013\22
Battlekat\Into the Forest (Dreamtrak Diamond Sound Remix)\2011\2013\23
Xeno & Oaklander\Sheen\2013\2013\24
Black Marble\A Great Design\2012\2013\25
Hypnotic School\Time for a Move (Steve Remix)\2013\2013\26
Douglas J. McCarthy\The Last Time\2012\2013\27
Blacksmif\...And the Sun Rose Out\2012\2013\28
Arnold Steiner\The Thinker\2013\2013\29
Chrissy Murderbot\Fuzzy\2012\2013\30
Nouvelle Phénomène\Au fond de mon coeur\2012\2013\31
Chvrches\ZVVL\2013\2013\32
Light Asylum\A Certain Person\2010\2013\33
Saint Etienne\Tonight\2012\2013\34
Molly Nilsson\I Hope You Die\2011\2013\35
Kobol Electronics\Dynatron\2011\2013\36
Jimmy Edgar\I Wanna be Your STD\2004\2013\37
Trust\The Last Dregs\2012\2013\38
Sally Shapiro\Lives Together\2013\2013\39
Rocket Lieber\Throw a Fit (DJ Clap Remix)\2011\2013\40
Boris Divider\Take My Beat\2004\2013\41
Pet Shop Boys\Inside a Dream\2013\2013\42
Clams Casino\Motivation\2011\2013\43
Kris Wadsworth\It's Time (Jimmy Edgar Remix)\2013\2013\44
Photodementia\Boxcia\2013\2013\45
Photodementia\Postpre\2013\2013\46
Machinedrum\Don't 1 2 Lose You\2013\2013\47
Kings of the Universe\Watching Over You\2012\2013\48
Bloom\Quartz (Starkey Remix)\2012\2013\49
Black Marble\Static\2012\2013\50
Disclosure\Lividup\2012\2013\51
Machinedrum\Gunshotta\2013\2013\52
Molly Nilsson\Dear Life\2013\2013\53
Brassica\At Least I Know Why\2013\2013\54
Hugh Masekela\Don't Go Lose it Baby (Stretch Mix)\1984\2013\55
Love You Long Time\I Had You Wrong (Kings of the Universe Remix)\2009\2013\56
Legowelt\Visions in My Mind\2013\2013\57
Plant43\Wounding Words\2012\2013\58
Trust\Shoom\2012\2013\59
Molly Nilsson\You Always Hurt the One You Love\2011\2013\60
Chvrches\Recover (Cid Rim Remix)\2013\2013\61
Bloom\Quartz (Slackk Remix)\2012\2013\62
Trust\F.T.F\2012\2013\63
EOD\Questionmark 3\2012\2013\64
Ortrotasce\World Unrelated\2013\2013\65
En Suite Cabinet\In Times (Version II)\2006\2013\66
Uexkull\Keonigs Division\2013\2013\67
Chvrches\Lies\2013\2013\68
Rene Bandaly Family\Tanki Tanki (Rabih Beaini Edit)\2012\2013\69
Molly Nilsson\City of Atlantis\2011\2013\70
Tangerine Dream\Hunting for Illusions\2011\2013\71
EOD\Arrow\2013\2013\72
Greystates\The Cult Of Mars\2012\2013\73
Exzakt\Clarity (Lethal Agent Remix)\2011\2013\74
Die Selektion\Gottes Wille\2013\2013\75
Parade Ground\Gold Rush\1987\2013\76
Niels Jensen\Propaganda\1984\2013\77
Dean Blunt and Inga Copeland\5\2012\2013\78
Sem\Red Dragon\1996\2013\79
Disclosure\Boiling\2012\2013\80
Saint Etienne\Over the Border\2012\2013\81
Photodementia\Synovium\2011\2013\82
Jean-Luc Ponty\In the Fast Lane\1989\2013\83
Black Marble\A Different Arrangement\2012\2013\84
Daniel Avery\Reception\2012\2013\85
Pet Shop Boys\Axis\2013\2013\86
Saint Etienne\Heading for the Fair\2012\2013\87
Cassie\King of Hearts (Richard X Remix)\2012\2013\88
Salma Agha\Come Closer\1984\2013\89
E.R.P.\Tuga\2013\2013\90
Pet Shop Boys\Vocal\2013\2013\91
Saint Etienne\I've Got Your Music\2012\2013\92
Ital Tek\Discontinuum\2012\2013\93
Molly Nilsson\Hotel Home\2011\2013\94
EOD\Innsmouth\2013\2013\95
Black Marble\MSQ No-Extra\2012\2013\96
Black Marble\UK\2012\2013\97
Scan 7\Black Moon Rising\1993\2013\98
Pet Shop Boys\Invisible\2012\2013\99
Pip Williams\Pressure Point\2011\2013\100
Machinedrum\The Statue\2011\2012\1
John Maus\This is the Beat\2005\2012\2
Blondes\Water (Bicep Remix)\2012\2012\3
John Maus\Castles in the Grave\2010\2012\4
Machinedrum\Now U Know Tha Deal 4 Real\2011\2012\5
Die Selektion\Raben\2011\2012\6
Vince Watson\Reach for the Sun\2012\2012\7
Trust\Sulk\2012\2012\8
Kuedo\Salt Lake Cuts\2011\2012\9
John Maus\Rights for Gays\2007\2012\10
TBA\The face we choose to miss\2011\2012\11
Kuedo\Work, Live & Sleep in Collapsing Space (Claude Speed 'Infinity Ultra Rework' feat. Jivraj Singh)\2012\2012\12
Die Selektion\Du rennst\2011\2012\13
The Shortwave Mystery\Signals from Afar (Vocalize)\1984\2012\14
Squarepusher\4001\2012\2012\15
Africa HiTech\Out in the Streets\2011\2012\16
Die Selektion\Deine Augen\2011\2012\17
Jessie Ware\Running (Disclosure Remix)\2012\2012\18
Kuedo\Vectoral\2011\2012\19
Eprom\Twerkul8\2011\2012\20
Salaligan\Samen\1983\2012\21
Current Value\Faith\2007\2012\22
B-Key\Man of Science\2011\2012\23
Logistics\Slow Motion\2008\2012\24
Squarepusher\Dark Steering\2012\2012\25
Björk\Thunderbolt (Current Value Remix)\2012\2012\26
Machinedrum\GBYE\2011\2012\27
Clio\Eyes (Extended Vocal Mix)\1984\2012\28
Squarepusher\Angel Integer\2012\2012\29
Die Selektion\Muskelberg (Kaleid Remix)\2011\2012\30
Grimes\Be a Body\2012\2012\31
Raiders of the Lost Arp\Lunar Lander\2011\2012\32
College feat. Electric Youth\A Real Hero\2009\2012\33
John Maus\Bennington\2007\2012\34
Sailor & I\Tough Love (Aril Brikha Remix)\2012\2012\35
Boris Divider\Citydrome\2012\2012\36
Mathew Jonson\Never Say Die (Remix)\2010\2012\37
Prurient\Palm Tree Corpse\2011\2012\38
Sunjammer\I Understand Now\2012\2012\39
John Maus\Don't Worship the Devil\2007\2012\40
Footprintz\Fear of Numbers\2012\2012\41
Son of Kick\Playing the Villain (Machinedrum Remix)\2011\2012\42
Led Er Est\Kaiyo Maru\2012\2012\43
Plant43\Fluid Reasoning\2012\2012\44
Kuedo\Ascension Phase\2011\2012\45
Kyau & Albert\Falling Anywhere (Sunn Jellie Remix)\2012\2012\46
Ital Tek\Pixel Haze\2012\2012\47
Ekman\Tears of a Clown (Video Version)\2012\2012\48
Distal\Behold The Jungle Bootleg\2012\2012\49
Timo Juuti & Hector 87\Cheap Bad Moves\2012\2012\50
Datassette\Partita for Unattended Computer\2012\2012\51
Vatican Shadow\September Cell (The Punishment)\2012\2012\52
Squarepusher\Energy Wizard\2012\2012\53
Björk\Solstice (Current Value Remix)\2012\2012\54
Tranzident & Peter Dubs\Drift (Daniel Kandi & Mark Andrez Rushed Mix)\2007\2012\55
B-Key\Uprising\2003\2012\56
Nu:Tone feat. Pat Fulgoni\Beliefs\2007\2012\57
Technicolour & Komatic\We Were Always One\2012\2012\58
Benoit & Sergio\Let Me Count the Ways (Extended Version)\2011\2012\59
Brassica\Made Up My Mind\2010\2012\60
Austra\The Villain\2011\2012\61
The Soul Drifters\Funky Soul Brother\1974\2012\62
Brassica\Lydden Circuit\2011\2012\63
Footprintz\Dangers Of the Mouth (Jimmy Edgar Remix)\2012\2012\64
Boris Divider\I Was\2012\2012\65
Vatican Shadow\Cairo is a Haunted City\2012\2012\66
Kuedo\Seeing the Edges\2011\2012\67
Ital Tek\Human Version\2012\2012\68
Dzeltenie Pastnieki\Kāpēc tu mani negribi\1982\2012\69
Die Selektion\Kühle Lippen\2011\2012\70
Die Selektion\Steine auf dein Haupt\2011\2012\71
John Maus\Too Much Money\2007\2012\72
Burial\Kindred\2012\2012\73
Claro Intelecto\Section (Part 2)\2004\2012\74
Austra\Beat and the Pulse\2010\2012\75
Donny & Current Value\Drill\2009\2012\76
Laurel Halo\Hour Logic\2011\2012\77
Conforce\24 (Gesloten Cirkel Remix)\2012\2012\78
Art Department\Tell Me Why (Part I)\2011\2012\79
Asha Puthli\Space Talk\1976\2012\80
Cause 4 Concern\Makes Me Wonder\2011\2012\81
Boris Divider\1983\2012\2012\82
Secret Squirrel\Jungle Squirrel (Juke Edit)\2011\2012\83
Machinedrum\Come1\2011\2012\84
Paradis\La Ballade de Jim\2011\2012\85
Dream Continuum\Giv a Lil Luv\2012\2012\86
xxxy\Ordinary Things\2011\2012\87
Dance Conspiracy\Dub War (Chapter Five)\1992\2012\88
Connan Mockasin\Forever Dolphin Love (Erol Alkan Rework)\2011\2012\89
Trust\Dressed for Space\2012\2012\90
Raiders of the Lost Arp\Night Theme\2011\2012\91
Paradis\Parfait Tirage\2011\2012\92
Legowelt\A Cold Winters Day\2012\2012\93
Martial Canterel\No Contact\2012\2012\94
Datassette\People Without Mouths\2012\2012\95
Jeremy Glenn\New Life (Perseus 'Summer of 83' Remix)\2011\2012\96
Fliehende Stürme\Stahl\2011\2012\97
DJ Taktix\Hornz For 94 (Philip D. Kick Footwork Edit)\2011\2012\98
Vince Watson\Found What I'm Looking for\2012\2012\99
Loreen\Euphoria\2012\2012\100
Emeli Sandé\Heaven\2011\2011\1
Pional\Into a Trap\2011\2011\2
Martial Canterel\Windscreen\2008\2011\3
John Maus\Head for the Country\2011\2011\4
The Dreams\Aloha Miami\2011\2011\5
John Maus\Streetlight\2011\2011\6
Det vackra livet\Viljan\2011\2011\7
Emeli Sandé\Heaven (Nu:Tone Remix)\2011\2011\8
Francisco\Moonroller (Raiders of the Lost Arp Mix)\2004\2011\9
Belong\Perfect Life\2011\2011\10
Martial Canterel\You Today\2010\2011\11
EOD\On a Herald Go\2010\2011\12
Datassette\Micro\2009\2011\13
Koreless\4D\2011\2011\14
Martial Canterel\Occupy These Terms\2011\2011\15
Vince Watson\My Desire\2009\2011\16
Vince Watson\Qualia\2009\2011\17
Vince Watson\Love in F Minor (Intro Mix)\2010\2011\18
Datassette\Flechte\2006\2011\19
Fet et Moi\Paris is for Lovers\2009\2011\20
Zouk Machine\A Pa Je (Smacked Out Mix)\2010\2011\21
John Maus\Keep Pushing On\2011\2011\22
Crystal Castles\Baptism\2010\2011\23
Starcluster feat. Marc Almond\Smoke & Mirrors (Starcluster Alternative Version)\2008\2011\24
Astrolabe\Leave the Station (Pelifics Remix)\2009\2011\25
John Maus\...and the Rain\2011\2011\26
D'Eon\Too Late to Choose\2010\2011\27
Balam Acab\Apart\2011\2011\28
Det vackra livet\Kristallen\2011\2011\29
Woodkid\Iron\2011\2011\30
Octo Octa\I'm Trying\2011\2011\31
John Maus\Quantum Leap\2011\2011\32
Nu:Tone\The Feeling\2011\2011\33
Pelifics feat. Miss Plug Inn\Andiamo al mare stanotte\2011\2011\34
Belong\Come See\2011\2011\35
Pional\Where Eagles Dare\2011\2011\36
Roberto Auser & Alden Tyrell\Blondes & Brunettes (Aldens Club Mix)\2010\2011\37
Candido\Thousand Finger Man\1979\2011\38
Manolo\Night Rhythm\2011\2011\39
Martial Canterel\Still a Part\2011\2011\40
Kuedo\Flight Path\2011\2011\41
The O'Jays\Put Our Heads Together\1983\2011\42
Pyramids with Nadja\An Angel Was Heard to Cry Over the City of Rome\2009\2011\43
John Maus\The Crucifix\2011\2011\44
Crystal Castles\Suffocation\2010\2011\45
Tangerine Dream\Horns of Doom\1985\2011\46
Marco Passarani\Nova\2008\2011\47
Limewax & Current Value\Tempest\2011\2011\48
Xeno & Oaklander\Sets & Lights\2011\2011\49
EOD\Utrecht\2010\2011\50
Xeno & Oaklander\Open Walls\2011\2011\51
Nu:Tone\Shine In\2011\2011\52
Datassette\The Aviatrix\2009\2011\53
Ndesh\Miserere Dub\2011\2011\54
Biosphere\Kobresia\1997\2011\55
Katy B feat. Magnetic Man\Perfect Stranger\2011\2011\56
CRC\Vaskitsaherra (E.R.P. aka Convextion Remix)\2009\2011\57
Xeno & Oaklander\Celeste\2008\2011\58
Miss Plug Inn\Sweetheart\2007\2011\59
Brassica\New Jam City\2010\2011\60
Teengirl Fantasy\Cheaters\2010\2011\61
Katy B\Broken Record\2011\2011\62
Octave One\I Believe (Sandwell District Remix)\2011\2011\63
Equip\XXXO\1983\2011\64
Crystal Castles\Vietnam\2010\2011\65
Det vackra livet\Askan\2011\2011\66
Martial Canterel\Secret Stores\2011\2011\67
John Maus\Hey Moon\2011\2011\68
Dexter\Junofest\2010\2011\69
Carol Jiani\Hit n Run Lover\1981\2011\70
Mr. Pauli\Der Alte\2008\2011\71
Niki & the Dove\DJ, Ease My Mind\2011\2011\72
Karl X Johan\Flames\2010\2011\73
Maja\If You Love Me Tonight (Passarani Mix)\2008\2011\74
D'Eon\Tear Down the Walls\2009\2011\75
Current Value\The Good\2009\2011\76
Space\Carry On Turn Me On\1977\2011\77
Martial Canterel\Some Days\2011\2011\78
Crystal Castles\Celestica\2010\2011\79
Det vackra livet\Barn av en istid\2011\2011\80
Gay Marvine\I'm Yr Money\2009\2011\81
Jules Tropicana\Come On\1983\2011\82
Maurice McGee\Do I Do\1983\2011\83
Danny Byrd\Shock Out\2008\2011\84
Totally Enormous Extinct Dinosaurs\Garden\2010\2011\85
Xeno & Oaklander\Italy\2011\2011\86
Xeno & Oaklander\Corrupt\2011\2011\87
Datashat\DCI Burnside\2011\2011\88
Dead Can Dance\How Fortunate the Man With None\1993\2011\89
Black Boned Angel\Verdun\2009\2011\90
Det vackra livet\Prärie av ljus\2011\2011\91
Elektridas\Elektridas\2009\2011\92
Professor Genius\Assassins (Time of the Assassins Steve Moore Remix)\2011\2011\93
SBTRKT\Pharaohs\2011\2011\94
Todd Terje\Snooze 4 Love\2011\2011\95
Wolfram\Hold My Breath (Sally Shapiro Version)\2011\2011\96
John Rocca\I Want it to be Real (Farley Mix)\1984\2011\97
Datassette\Space Rubbish Theme\2011\2011\98
Mehrwert\Man müsste Klavier spielen können\1982\2011\99
Poeme Electronique\My Complicated Personality\1982\2011\100
Games\Midi Drift\2010\2010\1
Oneohtrix Point Never\Physical Memory\2009\2010\2
E.R.P.\Frozen Volatiles\2010\2010\3
Xeno & Oaklander\4th Wall\2009\2010\4
Led Er Est\Scissors\2009\2010\5
Xeno & Oaklander\Shadow World\2009\2010\6
Games\Strawberry Skies\2010\2010\7
Romina Cohn\The Night\2001\2010\8
Fear of Tigers\I Can Make the Pain Disappear\2009\2010\9
Airiel\Thinktank\2007\2010\10
A Place to Bury Strangers\I Lived My Life to Stand in The Shadow of Your Heart\2009\2010\11
Cassie\Official Girl (CFCF Remix)\2008\2010\12
Gimmicks\Visst är du kär\1976\2010\13
Led Er Est\Port Isabel\2009\2010\14
XIX\1111.\2010\2010\15
Zola Jesus\Night\2010\2010\16
Fennesz\Rivers of Sand\2004\2010\17
Void Vision\In 20 Years\2010\2010\18
The Exaltics\Reticulation Notes\2009\2010\19
Xeno & Oaklander\Sentinelle\2009\2010\20
The Caretaker\Friends Past Re-United\2001\2010\21
Led Er Est\Laredo\2009\2010\22
Washed Out\Olivia\2009\2010\23
Xeno & Oaklander\Rendez-vous d'or\2009\2010\24
Sixfoe\Seasons\2004\2010\25
E.R.P.\El Camino\2010\2010\26
Oneohtrix Point Never\Betrayed in the Octagon\2007\2010\27
Ganymed\We Like You (The Way You Like Us)\1979\2010\28
Miss Kittin & The Hacker\1000 Dreams\2009\2010\29
Zola Jesus\Stridulum\2010\2010\30
Washed Out\Belong\2009\2010\31
Crystal Castles\Not in Love\2010\2010\32
Edrupt\M-U-S-I-K\2010\2010\33
Hurts\Wonderful Life\2010\2010\34
Washed Out\You'll See it\2009\2010\35
Liminals\The Swim\2009\2010\36
Xeno & Oaklander\Werke\2009\2010\37
oOoOO\Nosummr4U\2010\2010\38
Petit Mal\Song to Shout in the Ruins\2009\2010\39
Tiger & Woods\Gin Nation\2009\2010\40
Max & Intro\Beogradska Devojka\1984\2010\41
SSQ\Walkman On\1983\2010\42
Tensnake\Coma Cat\2010\2010\43
Urban Tribe\Insolitology\2010\2010\44
Liminals\Shine\2009\2010\45
Shamantis\J. Biebz - U Smile 800% Slower\2010\2010\46
Small Black\Despicable Dogs (Washed Out Remix)\2010\2010\47
Putsch '79\Samasaval\2010\2010\48
CFCF\It Was Never Meant to be this Way (Games Remix)\2010\2010\49
Washed Out\New Theory\2009\2010\50
Joker\Digidesign\2009\2010\51
Hudson Mohawke\Overnight\2009\2010\52
Passions\Endless\2010\2010\53
Fear of Tigers\Sirkka\2009\2010\54
Xeno & Oaklander\Saracen\2009\2010\55
Washed Out\Lately\2009\2010\56
Games\Shadows in Bloom\2010\2010\57
Disco Nihilist\Easy\2010\2010\58
Zola Jesus\Manifest Destiny\2010\2010\59
Linear Movement\Way Out of Living\1983\2010\60
Balam Acab\See Birds, Moon\2010\2010\61
Xeno & Oaklander\Preuss\2009\2010\62
Washed Out\Hold Out\2009\2010\63
Florence and the Machine\Rabbit Heart (Raise it Up) (Leo Zero Remix)\2009\2010\64
Hercules & Love Affair\You Belong\2008\2010\65
Oneohtrix Point Never\Zones Without People\2009\2010\66
Nocera\Let's go\1987\2010\67
Nadja\The Sun Always Shines on TV\2009\2010\68
The Mary Onettes\Void\2007\2010\69
Twisted Wires\Oh Hell\2010\2010\70
Led Er Est\The Unkept Area\2009\2010\71
Asso\Don't Stop\1983\2010\72
Oni Ayhun\OAR003-B\2009\2010\73
Ndesh\Grimeton\2010\2010\74
Bloodygrave & Die Lust!\Schnee in der Küche\2010\2010\75
Rustie\Bad Science\2009\2010\76
Polarkreis 18\Allein Allein\2008\2010\77
Azari & III\Hungry for the Power\2010\2010\78
Liars\Scissor\2009\2010\79
Enema & Gejonte\Mot nya djärva äventyr\1992\2010\80
Château Flight\Baltringue\2006\2010\81
Fear of Tigers\Calling Your Name\2009\2010\82
Lama\Nineteen Ninety Three\1983\2010\83
Salem\King Night\2010\2010\84
Grouper\Cover the Windows and the Walls\2007\2010\85
Julianna Barwick\Sunlight, Heaven\2009\2010\86
Enema & Gejonte\Mäklarnas dag\1992\2010\87
Gesloten Cirkel\Twisted Balloon\2009\2010\88
Belong\Same Places (Slow Version)\2008\2010\89
Liminals\Hands (for Rosemary Brown)\2009\2010\90
Rare Band\Why Why (Instrumental)\1986\2010\91
Xeno & Oaklander\Vagabond\2009\2010\92
Tensnake\Need Your Lovin\2010\2010\93
Balam Acab\Regret Making Mistakes\2010\2010\94
oOoOO\Burnout Eyess\2010\2010\95
Robin Thicke\Magic\2008\2010\96
Sophie Ellis-Bextor\Bittersweet\2010\2010\97
Oneohtrix Point Never\Hyperdawn\2008\2010\98
Nadja\Only Shallow\2009\2010\99
Underworld\Beautiful Burnout\2007\2010\100
Raiders of the Lost Arp\Azymuth\2008\2009\1
Hardfloor\The Trill Acid Theme (E.R.P. Remix)\2008\2009\2
Hardfloor\The Life We Choose (E.R.P. Remix)\2008\2009\3
Appaloosa\The Day (We Fell in Love)\2008\2009\4
House of House\Rushing to Paradise (Walkin' These Streets)\2009\2009\5
E.R.P.\Sensory Process\2009\2009\6
Guy Gerber\Timing\2009\2009\7
Moderat\Rusty Nails\2009\2009\8
Desire\If I Can't Hold You\2009\2009\9
Culoe De Song\The Bright Forest\2009\2009\10
Lykke Li\Breaking it Up (Familjen Remix)\2009\2009\11
Luomo\Love You All\2008\2009\12
College feat. Electric Youth\She Never Came Back (Russ Chimes Remix)\2008\2009\13
Barbara Morgenstern\Come to Berlin (Telefon Tel Aviv Mix)\2008\2009\14
52nd Street\Can't Afford\1984\2009\15
Bogdan Irkük a.k.a. Bulgari\Everything Is Changing\2008\2009\16
Telefon Tel Aviv\The Birds\2009\2009\17
Appaloosa\Intimate\2008\2009\18
Dosem\Beach Kisses (Rework)\2008\2009\19
Donna Summer\Now I Need You\1977\2009\20
Familjen\Det lilla livet\2007\2009\21
Hadamard\Spiritualisation of Cruelty\2007\2009\22
Gold Blood\She Doesn't Learn\2009\2009\23
Friday Bridge\This Case is Closed (Johan Agebjörn Remix)\2009\2009\24
Kings of the Universe\Acid Love\2009\2009\25
Spectrasoul\Alibi (Break Remix)\2009\2009\26
E.R.P.\Lodestone\2009\2009\27
Sally Shapiro\Let it Show\2009\2009\28
Appaloosa\Patchwork (Demo)\2008\2009\29
Mobius Band\The Loving Sounds of Static (Junior Boys Remix)\2006\2009\30
Hadamard\I Want to Know\2007\2009\31
Asobi Seksu\Me & Mary\2009\2009\32
Gold Blood\Another World\2009\2009\33
Abakus\Future Melt\2009\2009\34
Alisha\Baby Talk\1985\2009\35
Morgan Geist\24K\2001\2009\36
Friendly Fires feat. Au Revoir Simone\Paris (Aeroplane Remix)\2008\2009\37
Annie\Anthonio (Vaughn E Remix)\2009\2009\38
Gold Blood\On the Run\2009\2009\39
Pink Rhythm\Melodies of Love\1985\2009\40
Can\Future Days (Carl Craig Blade Runner Mix)\1997\2009\41
Klaus Schulze\Velvet Voyage\1977\2009\42
Koxo\Step by Step\1982\2009\43
Moreno\I Want to be Your Love Today\1986\2009\44
Manfred Mann\Just for Me\1968\2009\45
Gatekeeper\Optimus Maximus\2009\2009\46
Kaos\Definition of Love\1989\2009\47
Ada feat. Raz Ohara\Lovestoned\2009\2009\48
Dupont\Unknown Airspace\2004\2009\49
Rude 66\Fishbait\2008\2009\50
Real To Reel\Love Me Like This (Floating Points Remix)\2009\2009\51
The Naked Hearts\Only for You (Home Video Remix)\2009\2009\52
Rude 66\No One Had a Clue\2008\2009\53
Gavin Russom\The Fusion Point\2009\2009\54
Keen K & Dorian E\Lost But Not Found\2007\2009\55
Ronnie Dyson\All Over Your Face\1983\2009\56
David Joseph\You Can't Hide (Your Love From Me)\1983\2009\57
Moderat\Seamonkey\2009\2009\58
Bogdan Irkük a.k.a. Bulgari\Space Reflecting on the Bosporos\2008\2009\59
$tinkworx\Coelacanth\2008\2009\60
Motiivi:Tuntematon\1939\2005\2009\61
Sally Shapiro\Miracle\2009\2009\62
The Supremes\Let Yourself Go\1976\2009\63
Spewis\First and Last\2009\2009\64
Mount Kimbie\Maybes\2009\2009\65
Hieroglyphic Being\A Time Warp Synthesizer\2006\2009\66
Mathew Jonson\When Love Feels Like Crying\2009\2009\67
Motiivi:Tuntematon\I don't Feel Good (When You're not Around)\2007\2009\68
Sally Shapiro\Looking at the Stars\2009\2009\69
Morgan Geist\The Shore\2008\2009\70
Bat for Lashes\Daniel\2009\2009\71
Gold Blood\Well City\2009\2009\72
Box Codax\Missed Her Kiss\2006\2009\73
Brassica\Ballo dei Morti\2009\2009\74
The Juan Maclean\Happy House\2008\2009\75
Datassette\Weather Conditions\2009\2009\76
Beni\My Love Sees You (Classixx Remix)\2009\2009\77
Memory Cassette\Asleep at a Party\2009\2009\78
Melody Boy 2000\Monotone Fantastique (Monotone Mix)\1994\2009\79
Aeroplane\Caramellas\2007\2009\80
Hud Mo\Ooops!\2008\2009\81
Larry Young's Fuel\Turn Off The Lights\1975\2009\82
Rude 66\Walked The Line\2008\2009\83
Lime\You're My Magician\1981\2009\84
J.M. Silk\Shadows of Your Love (Ben Liebrand Minimix)\1986\2009\85
Erstlaub\Broadcasting on Ghost Frequencies (Part 1)\2009\2009\86
Meek Rabbit\Sweetheart in England\1984\2009\87
Kettel\Palle's Popsong\2008\2009\88
Lazer Crystal\Love Rhombus (Instrumental)\2009\2009\89
Kemal\Mutationz (Part 3)\2001\2009\90
Svreca\Eye (Hadamard Remix)\2009\2009\91
Kettel\The Wombat\2008\2009\92
Depeche Mode\Peace\2009\2009\93
Deadmau5 & Kaskade\I Remember\2008\2009\94
DJ Guy\Freak it All Night\2009\2009\95
Saint Etienne\Method of Modern Love (Cola Boy Mix)\2009\2009\96
Ndesh\Jetdaisuke FTW!!!\2009\2009\97
Cestrian\Mentor\2007\2009\98
Kris Menace presents Fred Falke\Fairlight\2006\2009\99
Xeno & Oaklander\Cold Forever\2007\2009\100
Jens Lekman\Sipping on the Sweet Nectar (Bogdan Irkük's Love Nectar Mix)\2008\2008\1
E.R.P.\Vox Automaton\2007\2008\2
Familjen\Huvudet i sanden\2007\2008\3
The Whitest Boy Alive\Golden Cage (Fred Falke Remix)\2008\2008\4
Tobiah\I Don't Really Exist\2006\2008\5
Tobiah\I Love Your Music\2006\2008\6
Fliehende Stürme\Lunaire\2008\2008\7
Slagsmålsklubben\Sponsored by Destiny\2007\2008\8
Tuxedomoon\In a Manner of Speaking\1985\2008\9
Cloetta Paris\Did We Collide?\2008\2008\10
Fall Of Saigon\She Leaves Me All Alone\1983\2008\11
Glass Candy\Life after Sundown\2007\2008\12
E.R.P.\Lament Subrosa\2007\2008\13
Lime\Babe, We're Gonna Love Tonight\1982\2008\14
Maximilian Skiba\Apple of Disco.Rd\2006\2008\15
Orgue Electronique\Die Liebe ist die größte Kraft\2005\2008\16
Maximilian Skiba\Violet Carnation\2006\2008\17
Starcluster feat. Elke B.\Jusqu'à la fin\2008\2008\18
Heartbreak\Akin to Dancing\2008\2008\19
Fixmer/McCarthy\Banging Down Your Door\2008\2008\20
Kleerup\Tower of Trellick\2008\2008\21
Mr. Clavio\Keine Gnade für die Sechste\2005\2008\22
Jesu\Friends are Evil\2004\2008\23
Kleerup feat. Neneh Cherry\Forever\2008\2008\24
Backlash\Lodestar\2006\2008\25
Asobi Seksu\Red Sea\2007\2008\26
Arvid Tuba\The Seasons are Sitting on Chairs\1998\2008\27
Vanessa van Basten\Floaters\2006\2008\28
Glass Domain\Interlock\1991\2008\29
Vanessa van Basten\Dole\2006\2008\30
Hjarnidaudi\March\2006\2008\31
Clashing Egos\Aminjig Nebere (I Trusted You) (Joakim's Afrobot mix)\2004\2008\32
Tracey Thorn\King's Cross (Hot Chip Remix)\2007\2008\33
Pride and Fall\Retrospect\2006\2008\34
Dream Disco\Take Me Home\2007\2008\35
Theo Parrish feat. Alena Waters\Soul Control\2007\2008\36
Frank Bolero\klkon\2007\2008\37
Quazar\The Seven Stars\1990\2008\38
Nu NRG\Bonsai\2004\2008\39
Pink Turns Blue\I Coldly Stare Out\1987\2008\40
Fliehende Stürme\Tobende Welt\2008\2008\41
Victrola\Maritime Tatami\1983\2008\42
Sally Shapiro\Jackie Jackie (Spend this Winter with Me) (Dyylan's Subzero Nocturne)\2008\2008\43
Oasis\Oasis Thirteen\2004\2008\44
Fliehende Stürme\Zuflucht\2008\2008\45
Pride and Fall\Border\2006\2008\46
Asobi Seksu\Thursday\2007\2008\47
Diode\No Mans Land\2007\2008\48
Fliehende Stürme\Kleines Herz\1999\2008\49
Forss\Journeyman\2003\2008\50
G.A.N.G.\KKK (Club Mix)\1983\2007\1
The Hasbeens\Make the World Go Away\2006\2007\2
Sally Shapiro\Skating in the Moonshine\2007\2007\3
Squadra Blanco\The Night Must Fall\2002\2007\4
Sally Shapiro\My Fantasy\2008\2007\5
Man Friday\Winners (Larry Levan Demo Mix)\1986\2007\6
Angie Care\Your Mind\1984\2007\7
Para One\Ski Lesson Blues\2006\2007\8
Legowelt\Congo Zombie\2005\2007\9
Rupesh Cartel\Ghost White (Ralf and Iza Remix)\2007\2007\10
Squarepusher\Planetarium\2006\2007\11
Above & Beyond\Alone Tonight\2006\2007\12
EMAK\Tanz in den Himmel\1982\2007\13
Sophie Rimheden feat. Annika Holmberg\Can You Save Me? (Mont Ventoux Remix)\2007\2007\14
Joe Yellow\Lover to Lover\1983\2007\15
Alba\Only Music Survives\1985\2007\16
Red White Rose\No one Puts Baby in the Corner\2003\2007\17
Din stalker\Herr Reporter\2007\2007\18
Legowelt\Hazy City Nights\2004\2007\19
Triola\Leuchtturm (Wighnomys Polarzip)\2005\2007\20
Komatrohn\Statist 2.0\2005\2007\21
Venise\Roissy\1988\2007\22
Sally Shapiro\Jackie Jackie (Spend this Winter with Me) (Dyylan's Subzero Nocturne)\2008\2007\23
Blank & Jones\Perfect Silence (Martin Roth Hardtrance Remix)\2004\2007\24
Zombi\Sapphire\2006\2007\25
Bloc Party\Where is Home? (Burial Remix)\2007\2007\26
Popular Computer\Next Level Pope\2006\2007\27
Covenant\The Men\2006\2007\28
Decadance\On and On (Fears Keep On) (Dub Version)\1983\2007\29
Thanya\Freedom\1982\2007\30
Den Harrow\Future Brain\1985\2007\31
Squarepusher\Tommib Help Buss\2004\2007\32
Kleerup feat. Robyn\With Every Heartbeat\2007\2007\33
Miss Kittin & The Hacker\Hometown\2007\2007\34
Sophie\Broken Tale\1986\2007\35
Annie\Heartbeat\2004\2007\36
Klapto\Mister Game (Alden Tyrell Vocal Remix)\2006\2007\37
Burial\Distant Lights\2006\2007\38
Ryuichi Sakamoto\The End Of Europe\1981\2007\39
Time\Holding On to love\1986\2007\40
DC Pöbeln med Guggi & 17\Bettan står i baren, baren är mitt mål, Bettan är baren\1985\2007\41
Simian Mobile Disco\It's the Beat (The Teenagers Remix)\2007\2007\42
Clio\Faces\1985\2007\43
Dennis Parker\Like an Eagle\1979\2007\44
Pascal F.E.O.S.\Synaptic\2006\2007\45
Change\The End\1980\2007\46
Heartbreak\We're Back\2007\2007\47
Cellophane\Music Colours\1984\2007\48
Johan Agebjörn\Mega Man II Re-mix\2007\2007\49
Polarius\Fallin Snow\2003\2007\50
Mark Tower\You aren't Fall in Love\1983\2007\51
The Field\Over the Ice\2007\2007\52
Oppenheimer Analysis\The Devil's Dancers\1982\2007\53
The Unknown Soldier\Babylon's Gifts\2006\2007\54
Blotnik Brothers\Love Song\2007\2007\55
Katy Gray\Hold Me Tight\1985\2007\56
Proceed\Laut\2007\2007\57
Papa Dance\W 40 dni dookola swiata\1984\2007\58
Purple Flash\We can Make it (1984 Instrumental)\1984\2007\59
Glass Candy\Miss Broadway\2007\2007\60
Junesex\Fast Food Messiahs (Carl A. Finlow Mix)\2004\2007\61
Daniel Wang\All Flowers Must Fade\2007\2007\62
Trilogy\Not Love\1982\2007\63
Para One\Liege\2006\2007\64
Covenant\Ritual Noise\2006\2007\65
Mike Mareen\Dancing in the Dark (Galactica Remix)\1985\2007\66
Umo Vogue\Just My Love\1984\2007\67
Ferry Corsten\Kyoto\2004\2007\68
Rhythm Talk\Groovin' (Active Club)\1984\2007\69
O'Gar\Playback Fantasy\1983\2007\70
Para One\Midnight Swim\2006\2007\71
Discomania\Everybody Wants to be Me\2004\2007\72
Mr. White\The Sun Can't Compare\2006\2007\73
Angel City\I Won't Let You Down\2005\2007\74
Cloetta Paris\Broken Heart Tango\2007\2007\75
Paul Hartnoll\Patchwork Guilt\2007\2007\76
Smith n Hack\Falling Stars\2007\2007\77
The Teenagers\Homecoming\2007\2007\78
New Baccara\Fantasy Boy\1988\2007\79
Above & Beyond\Tri-State\2006\2007\80
L.E.B. Harmony\Feeling Love\1978\2007\81
Vince Watson\MidiSensual\2006\2007\82
Covenant\Brave New World\2006\2007\83
Klaxons\Magick (Simian Mobile Disco Remix)\2007\2007\84
Squarepusher\Welcome to Europe\2006\2007\85
Above & Beyond\Hope\2006\2007\86
Wanexa\The Man from Colours\1982\2007\87
Antena\Camino Del Sol (Joakim Remix)\2006\2007\88
Mikado\Romance\1982\2007\89
Fox the Fox\Precious Little Diamond\1984\2007\90
LCD Soundsystem\Someone Great\2007\2007\91
Enter Shikari\Stand Your Ground; This is Ancient Land\2007\2007\92
Coco Bill\Evita\1984\2007\93
Aril Brikha\Last One\2007\2007\94
Ivan\Fotonovela\1984\2007\95
Prism\The White Shadow\1980\2007\96
Glass Candy\Rolling Down the Hills (Spring Demo)\2007\2007\97
Air France\Karibien\2006\2007\98
DJ Hell\Hot On the Heels of Love (Dave Clarke Remix)\1994\2007\99
Kai Del Noi\The Dream (Club Mix)\2005\2007\100
B.W.H.\Stop\1983\2006\1
Sally Shapiro\Hold Me So Tight\2006\2006\2
Sally Shapiro\I Know\2006\2006\3
Pineapples\Come On Closer\1983\2006\4
M & G\When I Let You Down\1986\2006\5
The Creatures\Believe in Yourself (Special Remix)\1983\2006\6
Sally Shapiro\Time to Let Go\2006\2006\7
The Expansives\Life with You\1982\2006\8
Severed Heads\Dead Eyes Opened\1984\2006\9
The Knife\The Captain\2006\2006\10
I.M.S.\Dancing Therapy\1984\2006\11
D.Kay + Raw.full\Bowser\2003\2006\12
M.I.K.E.\Lost My Way\2006\2006\13
Mr. Pauli feat. Mariana\Satisfaction\2006\2006\14
Ural 13 Diktators\Dream World\2001\2006\15
Freescha\Church Music\2002\2006\16
Ali Renault\Victory Horn\2005\2006\17
Kerri Chandler & Monique Bingham\In the Morning (Raw Mix)\2006\2006\18
Hugg & Pepp\Pellefant\2005\2006\19
Thomas Bronzwaer\Shadow World\2006\2006\20
I.M.S.\An English '93\1983\2006\21
Sally Shapiro\I'll be by Your Side\2006\2006\22
Spetsnaz\Totalitär\2006\2006\23
Gladio\Slave of Rome\2003\2006\24
Gentle Touch\Speaking of Reasonable\2006\2006\25
Klute\Hell Hath No Fury\2005\2006\26
VNV Nation\Airships\2002\2006\27
Ali Renault\Valentine\2005\2006\28
D'Malicious\Alive\2004\2006\29
Loui$\Magic Dance\1985\2006\30
Mew\Special\2005\2006\31
Technasia feat. Joris Voorn\'88 (All in All)\2006\2006\32
Armin van Buuren feat. Jan Vayne\Serenity\2005\2006\33
Frank Tavaglione\Tumidanda\1984\2006\34
VNV Nation\Beloved\2002\2006\35
Casco\Cybernetic Love\1983\2006\36
Daft Punk\The Prime Time of Your Life (Para One Remix)\NaN\2006\37
Junior Boys\So this is Goodbye\2006\2006\38
Mr. Pauli\Lo Mas\2006\2006\39
Sophie Rimheden\Queen of the Night (Rom Bansisco Mix)\2006\2006\40
Dharma\Plastic Doll\1982\2006\41
Rude 66\Overkill\2005\2006\42
Lo-Fi-Fnk\Change Channel\2006\2006\43
Yellow Magic Orchestra\Rydeen\1980\2006\44
Above and Beyond feat. Zoë Johnston\No One On Earth\2004\2006\45
Cyber People\Polaris\1984\2006\46
Airbase\Magic Silence (Intro)\2002\2006\47
Maximilian Skiba\Randez-vous\2005\2006\48
Dido\Take My Hand\1999\2006\49
M.I.K.E.\Voices from the Inside\2006\2006\50
Marco Passarani\Criticize\2005\2005\1
Pendulum\Masochist\2004\2005\2
The Light Bulb Project\Joystick\2004\2005\3
Joris Voorn\Incident\2004\2005\4
The Reese Project\The Colour Of Love (Underground Resistance Club Mix)\1992\2005\5
DJ Fresh\Submarines (Pendulum Remix)\2004\2005\6
The Radio Dept.\This Past Week\2005\2005\7
Ural 13 Diktators\Victorious Night\2000\2005\8
Duracell\Space Harrier/Turrican (Live at Barden's Boudoir)\2005\2005\9
Cat5\Sexy\2005\2005\10
Useless\Red X (Cymbalistic Remix by Dima)\2001\2005\11
Petter\These Days (Chable's Those Days Mix)\2005\2005\12
Nathan Fake\Dinamo\2005\2005\13
Mathew Jonson\Marionette\2004\2005\14
VNV Nation\Distant (Rubicon II)\1999\2005\15
The MFA\Motherload\2004\2005\16
VNV Nation\Darkangel\1999\2005\17
Breakage\Prophecy\2005\2005\18
Sushi\One More Chance\2005\2005\19
AFX\PWSteal.Ldpinch.D\2005\2005\20
Joris Voorn\Rejected\2004\2005\21
Extrawelt\Soopertrack\2005\2005\22
Ultrasonic\High Energy\2005\2005\23
Joris Voorn\Listen\2005\2005\24
E'Voke\Arms of Loren\1996\2005\25
VNV Nation\Saviour\1999\2005\26
Joris Voorn\Shining\2004\2005\27
The Radio Dept.\Deliverance\2005\2005\28
C-Bank\Perfect\1987\2005\29
Ariel Pink's Haunted Graffiti\Gray Sunset\2000\2005\30
Slam\Bright Lights Fading (Slam Return to Mono Mix)\2005\2005\31
Ficta\Eli\2004\2005\32
t.A.T.u.\Loves Me Not\2005\2005\33
Planisphere\Teardrop\2002\2005\34
The Radio Dept.\We Would Fall Against the Tide\2002\2005\35
AFX\I'm Self Employed\2005\2005\36
Lucknow Pact\Youth is for the Old\2005\2005\37
Lucknow Pact\A Few Drinks, a Few Laughs\2005\2005\38
Form & Function\Wonderland\2004\2005\39
Junkie XL\Today\2006\2005\40
Britney Spears\Breathe On Me (Holden Vocal)\2004\2005\41
Unai\Oh You And I (Trentemøller Mix)\2005\2005\42
Nitzer Ebb\Murderous (Phil Kieran Remix)\2004\2005\43
Trentemøller\Rykketid\2005\2005\44
Johannes Heil\Step into the Light\2004\2005\45
Midnight Star\Midas Touch (Hell Interface Remix)\1999\2005\46
The Light Bulb Project\Shine\2004\2005\47
Baxendale\I Built this City (Justus Köhncke Mix)\2005\2005\48
Junior Boys\Last Exit\2004\2005\49
Gino Soccio\Remember\1982\2005\50
